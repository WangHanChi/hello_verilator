      module our;
         initial begin $display("Hello World"); $finish; end
      endmodule    
	//our模块的功能是显示“Hello World"